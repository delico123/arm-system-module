module Extend(
	input clk,
	input [23:0] Instr,
	input [1:0] ImmSrc,
	output reg [31:0] ExtImm
	);

	always @(negedge clk)
		case(ImmSrc)
			// 8-bit unsigned immediate for data-processing
			2'b00: ExtImm = {24'b0, Instr[7:0]};
			// 12-bit unsigned immediate for LDR/STR
			2'b01: ExtImm = {20'b0, Instr[11:0]};
			// 24-bit two's complement(24-bit signed immediate) multiplied by 4 for Branch
			2'b10: ExtImm = {{6{Instr[23]}}, Instr[23:0], 2'b00};
			default: ExtImm = 32'bx; // undefined
	endcase
endmodule